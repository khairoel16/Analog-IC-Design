magic
tech sky130A
magscale 1 2
timestamp 1729221910
<< psubdiff >>
rect -262 1129 -202 1163
rect 946 1129 1006 1163
rect -262 1102 -228 1129
rect 972 1102 1006 1129
rect -262 -28 -228 -2
rect 972 -28 1006 -2
rect -262 -62 -202 -28
rect 946 -62 1006 -28
<< psubdiffcont >>
rect -202 1129 946 1163
rect -262 -2 -228 1102
rect 972 -2 1006 1102
rect -202 -62 946 -28
<< poly >>
rect -134 1082 -68 1098
rect -134 1048 -118 1082
rect -84 1048 -68 1082
rect -134 1032 -68 1048
rect -116 1006 -86 1032
rect 286 1028 458 1094
rect 812 1082 878 1098
rect 812 1048 828 1082
rect 862 1048 878 1082
rect 812 1032 878 1048
rect 270 518 474 584
rect -133 54 -67 70
rect -133 20 -117 54
rect -83 20 -67 54
rect -133 4 -67 20
rect 286 8 458 74
rect 813 54 879 70
rect 813 20 829 54
rect 863 20 879 54
rect 813 4 879 20
<< polycont >>
rect -118 1048 -84 1082
rect 828 1048 862 1082
rect -117 20 -83 54
rect 829 20 863 54
<< locali >>
rect -262 1129 -202 1163
rect 946 1129 1006 1163
rect -262 1102 -228 1129
rect 972 1102 1006 1129
rect -162 1048 -118 1082
rect -84 1048 -40 1082
rect -162 1006 -128 1048
rect -76 1032 -40 1048
rect -74 1006 -40 1032
rect 784 1048 828 1082
rect 862 1048 906 1082
rect 784 1010 818 1048
rect 870 1032 906 1048
rect 872 1010 906 1032
rect -162 70 -128 108
rect -74 70 -40 96
rect -162 54 -127 70
rect -75 54 -40 70
rect -162 20 -117 54
rect -83 20 -40 54
rect 782 54 819 108
rect 871 54 908 108
rect 782 20 829 54
rect 863 20 908 54
rect -262 -28 -228 -2
rect 972 -28 1006 -2
rect -262 -62 -202 -28
rect 946 -62 1006 -28
<< viali >>
rect 298 1129 332 1163
rect -118 1048 -84 1082
rect 828 1048 862 1082
rect -117 20 -83 54
rect 829 20 863 54
rect 412 -62 446 -28
<< metal1 >>
rect 286 1163 344 1169
rect 286 1129 298 1163
rect 332 1129 344 1163
rect -130 1082 -72 1088
rect -168 1048 -118 1082
rect -84 1081 -67 1082
rect -84 1048 -34 1081
rect -168 1042 -34 1048
rect -168 1006 -122 1042
rect -81 1032 -34 1042
rect -80 1006 -34 1032
rect 286 994 344 1129
rect 816 1082 874 1088
rect 778 1048 828 1082
rect 862 1081 879 1082
rect 862 1048 912 1081
rect 778 1042 912 1048
rect 778 1006 824 1042
rect 865 1032 912 1042
rect 866 1006 912 1032
rect -74 618 65 994
rect 279 690 289 994
rect 341 690 351 994
rect 393 618 403 994
rect 455 618 465 994
rect 624 618 634 994
rect 686 618 791 994
rect 31 606 65 618
rect 40 568 74 606
rect 40 534 704 568
rect 670 484 704 534
rect -74 108 2 484
rect 58 108 74 484
rect 279 108 289 484
rect 341 108 351 484
rect 393 108 403 412
rect 455 108 465 412
rect 670 108 818 484
rect -168 60 -122 108
rect -80 60 -34 108
rect -168 54 -34 60
rect -168 20 -117 54
rect -83 20 -34 54
rect -129 14 -71 20
rect 400 -28 458 108
rect 778 60 824 108
rect 866 60 912 108
rect 778 54 912 60
rect 778 20 829 54
rect 863 20 912 54
rect 817 14 875 20
rect 400 -62 412 -28
rect 446 -62 458 -28
rect 400 -68 458 -62
<< via1 >>
rect 289 690 341 994
rect 403 618 455 994
rect 634 618 686 994
rect 2 108 58 484
rect 289 108 341 484
rect 403 108 455 412
<< metal2 >>
rect 287 994 343 1004
rect 287 680 343 690
rect 403 994 455 1004
rect 403 572 455 618
rect 632 994 688 1004
rect 632 608 688 618
rect 289 530 455 572
rect 2 484 58 494
rect 2 98 58 108
rect 289 484 341 530
rect 289 98 341 108
rect 401 412 457 422
rect 401 98 457 108
<< via2 >>
rect 287 690 289 994
rect 289 690 341 994
rect 341 690 343 994
rect 632 618 634 994
rect 634 618 686 994
rect 686 618 688 994
rect 2 108 58 484
rect 401 108 403 412
rect 403 108 455 412
rect 455 108 457 412
<< metal3 >>
rect 277 994 353 999
rect 622 994 698 999
rect 273 690 283 994
rect 347 690 357 994
rect 277 685 353 690
rect 622 618 632 994
rect 688 618 698 994
rect 622 613 698 618
rect 622 580 690 613
rect -8 520 690 580
rect -8 484 68 520
rect -8 108 2 484
rect 58 108 68 484
rect 391 412 467 417
rect 387 108 397 412
rect 461 108 471 412
rect -8 103 68 108
rect 391 103 467 108
<< via3 >>
rect 283 690 287 994
rect 287 690 343 994
rect 343 690 347 994
rect 397 108 401 412
rect 401 108 457 412
rect 457 108 461 412
<< metal4 >>
rect 282 994 348 995
rect 282 690 283 994
rect 347 690 348 994
rect 273 585 357 690
rect 273 517 471 585
rect 387 412 471 517
rect 396 108 397 412
rect 461 108 462 412
rect 396 107 462 108
use sky130_fd_pr__nfet_01v8_4HFSKE  sky130_fd_pr__nfet_01v8_4HFSKE_0
timestamp 1729216608
transform 1 0 845 0 1 806
box -73 -226 73 226
use sky130_fd_pr__nfet_01v8_4HFSKE  sky130_fd_pr__nfet_01v8_4HFSKE_1
timestamp 1729216608
transform 1 0 -101 0 1 806
box -73 -226 73 226
use sky130_fd_pr__nfet_01v8_4HFSKE  sky130_fd_pr__nfet_01v8_4HFSKE_2
timestamp 1729216608
transform 1 0 -101 0 1 296
box -73 -226 73 226
use sky130_fd_pr__nfet_01v8_4HFSKE  sky130_fd_pr__nfet_01v8_4HFSKE_3
timestamp 1729216608
transform 1 0 845 0 1 296
box -73 -226 73 226
use sky130_fd_pr__nfet_01v8_QCS68M  sky130_fd_pr__nfet_01v8_QCS68M_0
timestamp 1729216608
transform 1 0 372 0 1 551
box -344 -543 344 543
<< labels >>
flabel space 153 812 161 817 0 FreeSans 320 0 0 0 M3
flabel via1 306 892 314 897 0 FreeSans 320 0 0 0 S3
flabel space 552 819 560 824 0 FreeSans 320 0 0 0 M4
flabel space 553 329 561 334 0 FreeSans 320 0 0 0 M3
flabel space 189 323 197 328 0 FreeSans 320 0 0 0 M4
flabel via1 310 394 318 399 0 FreeSans 320 0 0 0 S4
flabel via1 424 894 432 899 0 FreeSans 320 0 0 0 S4
flabel via1 426 405 434 410 0 FreeSans 320 0 0 0 S3
flabel via1 656 900 664 905 0 FreeSans 320 0 0 0 D4
flabel metal1 685 395 693 400 0 FreeSans 320 0 0 0 D3
flabel metal1 54 830 54 830 0 FreeSans 320 0 0 0 D3
flabel metal1 2 745 2 745 0 FreeSans 320 0 0 0 D3
port 1 nsew
flabel metal2 427 595 427 595 0 FreeSans 320 0 0 0 RS
port 2 nsew
flabel metal3 678 588 678 588 0 FreeSans 320 0 0 0 D4
port 4 nsew
flabel viali 431 -42 431 -42 0 FreeSans 320 0 0 0 GND
port 6 nsew
<< end >>
