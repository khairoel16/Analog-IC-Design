magic
tech sky130A
magscale 1 2
timestamp 1729323365
<< nwell >>
rect -297 -258 1402 1094
<< nsubdiff >>
rect -261 1024 -201 1058
rect 1306 1024 1366 1058
rect -261 994 -227 1024
rect 1332 994 1366 1024
rect -261 -188 -227 -166
rect 1332 -188 1366 -166
rect -261 -222 -201 -188
rect 1306 -222 1366 -188
<< nsubdiffcont >>
rect -201 1024 1306 1058
rect -261 -166 -227 994
rect 1332 -166 1366 994
rect -201 -222 1306 -188
<< poly >>
rect -126 838 -60 854
rect -126 804 -110 838
rect -76 804 -60 838
rect -126 788 -60 804
rect 1165 838 1231 854
rect 1165 804 1181 838
rect 1215 804 1231 838
rect 1165 788 1231 804
rect -108 762 -78 788
rect 1182 760 1212 788
rect -108 69 -78 75
rect 1182 69 1212 100
rect -125 53 -59 69
rect -125 19 -109 53
rect -75 19 -59 53
rect -125 3 -59 19
rect 1164 53 1230 69
rect 1164 19 1180 53
rect 1214 19 1230 53
rect 1164 3 1230 19
<< polycont >>
rect -110 804 -76 838
rect 1181 804 1215 838
rect -109 19 -75 53
rect 1180 19 1214 53
<< locali >>
rect -261 1024 -201 1058
rect 1306 1024 1366 1058
rect -261 994 -227 1024
rect 1332 994 1366 1024
rect -154 804 -110 838
rect -76 804 -32 838
rect -154 736 -120 804
rect -66 736 -32 804
rect 1136 804 1181 838
rect 1215 804 1258 838
rect 1136 740 1170 804
rect 1224 738 1258 804
rect -154 53 -120 97
rect -66 53 -32 98
rect -154 19 -109 53
rect -75 19 -32 53
rect 1136 53 1170 96
rect 1224 53 1258 96
rect 1136 19 1180 53
rect 1214 19 1258 53
rect -154 13 -120 19
rect -261 -188 -227 -166
rect 1332 -188 1366 -166
rect -261 -222 -201 -188
rect 1306 -222 1366 -188
<< viali >>
rect -110 804 -76 838
rect 1181 804 1215 838
rect -109 19 -75 53
rect 1180 19 1214 53
rect 518 -222 585 -188
<< metal1 >>
rect 218 855 886 883
rect -122 838 -64 844
rect -160 804 -110 838
rect -76 804 -26 838
rect -160 798 -26 804
rect -160 724 -114 798
rect -72 736 -26 798
rect -72 724 82 736
rect 218 724 246 855
rect 490 724 518 855
rect 586 724 614 855
rect 858 724 886 855
rect 1130 838 1264 844
rect 1130 804 1181 838
rect 1215 804 1264 838
rect 1130 798 1264 804
rect 1130 730 1176 798
rect 1218 730 1264 798
rect -66 670 82 724
rect 1022 670 1170 724
rect -66 607 39 670
rect 91 607 101 670
rect 301 607 311 670
rect 363 607 373 670
rect 731 607 741 670
rect 793 607 803 670
rect 1003 607 1013 670
rect 1065 607 1170 670
rect -66 548 82 607
rect 1022 548 1170 607
rect -72 536 82 548
rect -72 444 -26 536
rect 30 444 40 500
rect 100 446 110 498
rect 178 446 188 498
rect 372 446 382 498
rect 450 446 460 498
rect -226 336 -216 392
rect -160 336 -26 392
rect 100 338 110 390
rect 178 338 188 390
rect 372 338 382 390
rect 450 338 460 390
rect -72 293 -26 336
rect 490 288 518 548
rect 586 288 614 548
rect 1130 500 1176 539
rect 644 446 654 498
rect 722 446 732 498
rect 916 446 926 498
rect 994 446 1004 498
rect 1130 444 1264 500
rect 1320 444 1330 500
rect 644 338 654 390
rect 722 338 732 390
rect 916 338 926 390
rect 994 338 1004 390
rect 1064 336 1074 392
rect 1130 300 1176 392
rect -66 229 82 288
rect 1022 229 1170 288
rect -66 166 39 229
rect 91 166 101 229
rect 301 166 311 229
rect 363 166 373 229
rect 731 166 741 229
rect 793 166 803 229
rect 1003 166 1013 229
rect 1065 166 1170 229
rect -66 112 82 166
rect 1022 112 1170 166
rect -160 59 -114 101
rect -72 59 -26 106
rect -160 53 -26 59
rect -160 19 -109 53
rect -75 19 -26 53
rect -160 13 -63 19
rect 218 -37 246 112
rect 490 -37 518 112
rect 586 -37 614 112
rect 858 -37 886 112
rect 1130 59 1176 100
rect 1218 59 1264 100
rect 1130 53 1264 59
rect 1130 19 1180 53
rect 1214 19 1264 53
rect 1130 13 1264 19
rect 218 -65 886 -37
rect 506 -188 597 -182
rect 506 -222 518 -188
rect 585 -222 597 -188
rect 506 -228 597 -222
<< via1 >>
rect 39 607 91 670
rect 311 607 363 670
rect 741 607 793 670
rect 1013 607 1065 670
rect -26 444 30 500
rect 110 446 178 498
rect 382 446 450 498
rect -216 336 -160 392
rect 110 338 178 390
rect 382 338 450 390
rect 654 446 722 498
rect 926 446 994 498
rect 1264 444 1320 500
rect 654 338 722 390
rect 926 338 994 390
rect 1074 336 1130 392
rect 39 166 91 229
rect 311 166 363 229
rect 741 166 793 229
rect 1013 166 1065 229
<< metal2 >>
rect 39 855 363 907
rect 39 670 91 855
rect 39 597 91 607
rect 311 670 363 855
rect 311 597 363 607
rect 741 855 1065 907
rect 741 670 793 855
rect 741 597 793 607
rect 1013 670 1065 855
rect 1013 597 1065 607
rect -26 500 30 510
rect 450 508 586 509
rect -26 434 30 444
rect 110 498 586 508
rect 178 446 382 498
rect 450 446 586 498
rect 110 437 586 446
rect 110 436 450 437
rect -216 392 -160 402
rect -216 326 -160 336
rect 110 392 178 402
rect 110 326 178 336
rect 382 392 450 402
rect 382 326 450 336
rect 518 401 586 437
rect 654 500 722 510
rect 654 434 722 444
rect 926 500 994 510
rect 926 434 994 444
rect 1264 500 1320 510
rect 1264 434 1320 444
rect 518 400 722 401
rect 518 390 994 400
rect 518 338 654 390
rect 722 338 926 390
rect 518 328 994 338
rect 1074 392 1130 402
rect 1074 326 1130 336
rect 39 229 91 239
rect 39 -19 91 166
rect 311 229 363 239
rect 311 -19 363 166
rect 39 -71 363 -19
rect 741 229 793 239
rect 741 -19 793 166
rect 1013 229 1065 239
rect 1013 -19 1065 166
rect 741 -71 1065 -19
<< via2 >>
rect -26 444 30 500
rect -216 336 -160 392
rect 110 390 178 392
rect 110 338 178 390
rect 110 336 178 338
rect 382 390 450 392
rect 382 338 450 390
rect 382 336 450 338
rect 654 498 722 500
rect 654 446 722 498
rect 654 444 722 446
rect 926 498 994 500
rect 926 446 994 498
rect 926 444 994 446
rect 1264 444 1320 500
rect 1074 336 1130 392
<< metal3 >>
rect -226 956 1330 1018
rect -226 392 -150 956
rect -226 336 -216 392
rect -160 336 -150 392
rect -226 -120 -150 336
rect -36 833 1140 896
rect -36 500 40 833
rect -36 444 -26 500
rect 30 444 40 500
rect -36 3 40 444
rect 518 500 1004 505
rect 518 444 654 500
rect 722 444 926 500
rect 994 444 1004 500
rect 518 439 1004 444
rect 518 397 586 439
rect 100 392 586 397
rect 100 336 110 392
rect 178 336 382 392
rect 450 336 586 392
rect 100 331 586 336
rect 1064 392 1140 833
rect 1064 336 1074 392
rect 1130 336 1140 392
rect 1064 3 1140 336
rect -36 -60 1140 3
rect 1254 500 1330 956
rect 1254 444 1264 500
rect 1320 444 1330 500
rect 1254 -120 1330 444
rect -226 -182 1330 -120
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_0
timestamp 1729241875
transform 1 0 1197 0 1 636
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_1
timestamp 1729241875
transform 1 0 -93 0 1 200
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_2
timestamp 1729241875
transform 1 0 1197 0 1 200
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_3
timestamp 1729241875
transform 1 0 -93 0 1 636
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_FH5654  sky130_fd_pr__pfet_01v8_FH5654_0
timestamp 1729239931
transform 1 0 552 0 1 418
box -552 -418 552 418
<< labels >>
flabel nwell 414 651 420 652 0 FreeSans 160 0 0 0 M6
flabel nwell 688 201 694 202 0 FreeSans 160 0 0 0 M6
flabel nwell 689 641 695 642 0 FreeSans 160 0 0 0 M7
flabel nwell 414 194 420 195 0 FreeSans 160 0 0 0 M7
flabel nwell 148 201 154 202 0 FreeSans 160 0 0 0 M7
flabel via1 335 646 335 646 0 FreeSans 160 0 0 0 d6
flabel via1 63 646 63 646 0 FreeSans 160 0 0 0 d6
flabel via1 1036 196 1036 196 0 FreeSans 160 0 0 0 d6
flabel via1 768 198 768 198 0 FreeSans 160 0 0 0 d6
flabel nwell 964 646 970 647 0 FreeSans 160 0 0 0 M7
flabel nwell 962 200 968 201 0 FreeSans 160 0 0 0 M6
flabel nwell 140 648 146 649 0 FreeSans 160 0 0 0 M6
flabel nwell 550 -207 552 -206 0 FreeSans 160 0 0 0 VDD
port 8 nsew
flabel metal1 597 796 597 796 0 FreeSans 160 0 0 0 D5
port 13 nsew
flabel metal2 324 795 324 795 0 FreeSans 160 0 0 0 D6
port 22 nsew
flabel metal3 815 473 815 473 0 FreeSans 160 0 0 0 VIP
port 23 nsew
flabel via1 767 638 767 638 0 FreeSans 160 0 0 0 d7
flabel via1 331 201 331 201 0 FreeSans 160 0 0 0 d7
flabel metal2 331 53 331 53 0 FreeSans 160 0 0 0 OUT
port 26 nsew
flabel metal2 276 473 276 473 0 FreeSans 160 0 0 0 VIN
port 28 nsew
flabel via1 1043 649 1043 649 0 FreeSans 160 0 0 0 d7
<< end >>
