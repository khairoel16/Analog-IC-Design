magic
tech sky130A
magscale 1 2
timestamp 1729407323
<< nwell >>
rect -2443 2244 -1441 2650
rect -1499 320 -1444 510
rect -1499 316 -1442 320
rect -1499 -624 -1242 316
rect -2440 -628 -1242 -624
rect -2441 -823 -1242 -628
rect -2442 -859 423 -823
rect -2443 -866 423 -859
rect -2443 -1036 -1276 -866
<< metal1 >>
rect -1258 2228 -1212 2253
rect -1460 2164 -1450 2228
rect -1382 2164 -1212 2228
rect -1004 1755 -865 1790
rect -461 1622 -391 1634
rect -804 1573 162 1622
rect -1452 1436 -1216 1502
rect -1452 857 -1382 1436
rect 92 1085 162 1573
rect 328 1374 338 1515
rect 488 1374 498 1515
rect 328 1177 338 1318
rect 488 1177 498 1318
rect 328 1085 338 1120
rect 92 1015 338 1085
rect 328 979 338 1015
rect 488 979 498 1120
rect 328 889 338 923
rect -1790 851 -1382 857
rect -1850 795 -1840 851
rect -1784 795 -1382 851
rect -1790 788 -1382 795
rect 92 819 338 889
rect -1234 408 -1224 475
rect -1162 408 -1152 475
rect 92 336 162 819
rect 328 782 338 819
rect 488 782 498 923
rect 328 584 338 725
rect 488 584 498 725
rect 328 394 338 535
rect 488 394 498 535
rect 379 393 449 394
rect -473 287 162 336
rect -473 285 -382 287
rect -199 -446 -189 -382
rect -121 -446 -111 -382
rect -1850 -526 -1840 -459
rect -1778 -526 -1768 -459
rect -1628 -870 -1558 -479
rect -462 -870 -392 -812
rect -1628 -919 -392 -870
<< via1 >>
rect -1450 2164 -1382 2228
rect 338 1374 488 1515
rect 338 1177 488 1318
rect 338 979 488 1120
rect -1840 795 -1784 851
rect -1224 408 -1162 475
rect 338 782 488 923
rect 338 584 488 725
rect 338 394 488 535
rect -189 -446 -121 -382
rect -1840 -526 -1778 -459
<< metal2 >>
rect -1450 2228 -1382 2238
rect -1450 2154 -1382 2164
rect -736 1969 -668 1979
rect -736 1895 -668 1905
rect -695 1573 247 1622
rect -695 1394 -627 1573
rect 177 1280 247 1573
rect 338 1515 488 1525
rect 338 1364 488 1374
rect 338 1318 488 1328
rect 177 1210 338 1280
rect 338 1167 488 1177
rect 338 1120 488 1130
rect 338 969 488 979
rect 338 923 488 933
rect -1840 851 -1784 861
rect -1840 785 -1784 795
rect 338 772 488 782
rect 338 725 488 735
rect 177 623 338 693
rect -1224 476 -1162 485
rect -1452 475 -1162 476
rect -1452 408 -1224 475
rect -1452 407 -1162 408
rect -1840 -458 -1778 -449
rect -1452 -458 -1382 407
rect -1224 398 -1162 407
rect 177 337 247 623
rect 338 574 488 584
rect 338 535 488 545
rect 338 384 488 394
rect -461 286 247 337
rect -461 -273 -393 286
rect -189 -382 -121 -372
rect -189 -456 -121 -446
rect -1840 -459 -1382 -458
rect -1778 -526 -1382 -459
rect -1840 -527 -1382 -526
rect -1840 -536 -1778 -527
<< via2 >>
rect -1450 2164 -1382 2228
rect -736 1905 -668 1969
rect 338 1374 488 1515
rect -189 -446 -121 -382
<< metal3 >>
rect -1460 2228 -1372 2233
rect -1460 2164 -1450 2228
rect -1382 2164 -1372 2228
rect -1460 1669 -1372 2164
rect -746 1969 -658 1974
rect -746 1905 -736 1969
rect -668 1905 -658 1969
rect -746 1900 -658 1905
rect -736 1632 -668 1900
rect -736 1564 0 1632
rect -70 1478 0 1564
rect 328 1515 498 1520
rect 328 1478 338 1515
rect -70 1418 338 1478
rect -70 178 0 1418
rect 328 1374 338 1418
rect 488 1374 498 1515
rect 328 1369 498 1374
rect 328 394 338 535
rect 488 394 498 535
rect -1019 -445 -1009 -381
rect -941 -445 -931 -381
rect -199 -382 -111 -377
rect -199 -446 -189 -382
rect -121 -446 -111 -382
rect -199 -451 -111 -446
<< via3 >>
rect -1450 2164 -1382 2228
rect 338 394 488 535
rect -1009 -445 -941 -381
rect -189 -446 -121 -382
<< metal4 >>
rect -1460 2228 -1372 2229
rect -1460 2164 -1450 2228
rect -1382 2164 -1372 2228
rect -1460 -380 -1372 2164
rect 337 535 489 536
rect 337 494 338 535
rect 17 434 338 494
rect 17 346 77 434
rect 337 394 338 434
rect 488 394 489 535
rect 337 393 489 394
rect -190 286 77 346
rect -1460 -381 -940 -380
rect -1460 -417 -1009 -381
rect -1459 -445 -1009 -417
rect -941 -445 -940 -381
rect -1459 -446 -940 -445
rect -190 -382 -120 286
rect -190 -446 -189 -382
rect -121 -446 -120 -382
rect -190 -447 -120 -446
use nmoscs  nmoscs_0
timestamp 1729221910
transform 1 0 -1090 0 1 404
box -262 -68 1006 1169
use nmosds  nmosds_0
timestamp 1729235038
transform -1 0 210 0 -1 2533
box -290 -116 1562 910
use pmoscs2  pmoscs2_0
timestamp 1729323365
transform 1 0 -979 0 -1 58
box -297 -258 1402 1094
use pmoscs  pmoscs_0
timestamp 1729163496
transform 1 0 -2261 0 1 366
box -179 -1003 819 1915
<< labels >>
flabel metal3 395 1444 398 1444 0 FreeSans 480 0 0 0 OUT
port 1 nsew
flabel via1 414 1250 414 1250 0 FreeSans 480 0 0 0 RS
port 2 nsew
flabel via1 420 1040 420 1040 0 FreeSans 480 0 0 0 GND
port 3 nsew
flabel via1 406 843 406 843 0 FreeSans 480 0 0 0 VDD
port 4 nsew
flabel via1 403 654 403 654 0 FreeSans 480 0 0 0 VIN
port 5 nsew
flabel via3 409 458 409 458 0 FreeSans 480 0 0 0 VIP
port 7 nsew
<< end >>
