magic
tech sky130A
magscale 1 2
timestamp 1729224540
<< nmos >>
rect -407 47 -247 247
rect -189 47 -29 247
rect 29 47 189 247
rect 247 47 407 247
rect -407 -247 -247 -47
rect -189 -247 -29 -47
rect 29 -247 189 -47
rect 247 -247 407 -47
<< ndiff >>
rect -465 235 -407 247
rect -465 59 -453 235
rect -419 59 -407 235
rect -465 47 -407 59
rect -247 235 -189 247
rect -247 59 -235 235
rect -201 59 -189 235
rect -247 47 -189 59
rect -29 235 29 247
rect -29 59 -17 235
rect 17 59 29 235
rect -29 47 29 59
rect 189 235 247 247
rect 189 59 201 235
rect 235 59 247 235
rect 189 47 247 59
rect 407 235 465 247
rect 407 59 419 235
rect 453 59 465 235
rect 407 47 465 59
rect -465 -59 -407 -47
rect -465 -235 -453 -59
rect -419 -235 -407 -59
rect -465 -247 -407 -235
rect -247 -59 -189 -47
rect -247 -235 -235 -59
rect -201 -235 -189 -59
rect -247 -247 -189 -235
rect -29 -59 29 -47
rect -29 -235 -17 -59
rect 17 -235 29 -59
rect -29 -247 29 -235
rect 189 -59 247 -47
rect 189 -235 201 -59
rect 235 -235 247 -59
rect 189 -247 247 -235
rect 407 -59 465 -47
rect 407 -235 419 -59
rect 453 -235 465 -59
rect 407 -247 465 -235
<< ndiffc >>
rect -453 59 -419 235
rect -235 59 -201 235
rect -17 59 17 235
rect 201 59 235 235
rect 419 59 453 235
rect -453 -235 -419 -59
rect -235 -235 -201 -59
rect -17 -235 17 -59
rect 201 -235 235 -59
rect 419 -235 453 -59
<< poly >>
rect -407 247 -247 273
rect -189 247 -29 273
rect 29 247 189 273
rect 247 247 407 273
rect -407 21 -247 47
rect -189 21 -29 47
rect 29 21 189 47
rect 247 21 407 47
rect -407 -47 -247 -21
rect -189 -47 -29 -21
rect 29 -47 189 -21
rect 247 -47 407 -21
rect -407 -273 -247 -247
rect -189 -273 -29 -247
rect 29 -273 189 -247
rect 247 -273 407 -247
<< locali >>
rect -453 235 -419 251
rect -453 43 -419 59
rect -235 235 -201 251
rect -235 43 -201 59
rect -17 235 17 251
rect -17 43 17 59
rect 201 235 235 251
rect 201 43 235 59
rect 419 235 453 251
rect 419 43 453 59
rect -453 -59 -419 -43
rect -453 -251 -419 -235
rect -235 -59 -201 -43
rect -235 -251 -201 -235
rect -17 -59 17 -43
rect -17 -251 17 -235
rect 201 -59 235 -43
rect 201 -251 235 -235
rect 419 -59 453 -43
rect 419 -251 453 -235
<< viali >>
rect -453 59 -419 235
rect -235 59 -201 235
rect -17 59 17 235
rect 201 59 235 235
rect 419 59 453 235
rect -453 -235 -419 -59
rect -235 -235 -201 -59
rect -17 -235 17 -59
rect 201 -235 235 -59
rect 419 -235 453 -59
<< metal1 >>
rect -459 235 -413 247
rect -459 59 -453 235
rect -419 59 -413 235
rect -459 47 -413 59
rect -241 235 -195 247
rect -241 59 -235 235
rect -201 59 -195 235
rect -241 47 -195 59
rect -23 235 23 247
rect -23 59 -17 235
rect 17 59 23 235
rect -23 47 23 59
rect 195 235 241 247
rect 195 59 201 235
rect 235 59 241 235
rect 195 47 241 59
rect 413 235 459 247
rect 413 59 419 235
rect 453 59 459 235
rect 413 47 459 59
rect -459 -59 -413 -47
rect -459 -235 -453 -59
rect -419 -235 -413 -59
rect -459 -247 -413 -235
rect -241 -59 -195 -47
rect -241 -235 -235 -59
rect -201 -235 -195 -59
rect -241 -247 -195 -235
rect -23 -59 23 -47
rect -23 -235 -17 -59
rect 17 -235 23 -59
rect -23 -247 23 -235
rect 195 -59 241 -47
rect 195 -235 201 -59
rect 235 -235 241 -59
rect 195 -247 241 -235
rect 413 -59 459 -47
rect 413 -235 419 -59
rect 453 -235 459 -59
rect 413 -247 459 -235
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1 l 0.8 m 2 nf 4 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 70 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
