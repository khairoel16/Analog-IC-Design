magic
tech sky130A
magscale 1 2
timestamp 1729224540
<< nmos >>
rect -407 109 -247 309
rect -189 109 -29 309
rect 29 109 189 309
rect 247 109 407 309
rect -407 -309 -247 -109
rect -189 -309 -29 -109
rect 29 -309 189 -109
rect 247 -309 407 -109
<< ndiff >>
rect -465 297 -407 309
rect -465 121 -453 297
rect -419 121 -407 297
rect -465 109 -407 121
rect -247 297 -189 309
rect -247 121 -235 297
rect -201 121 -189 297
rect -247 109 -189 121
rect -29 297 29 309
rect -29 121 -17 297
rect 17 121 29 297
rect -29 109 29 121
rect 189 297 247 309
rect 189 121 201 297
rect 235 121 247 297
rect 189 109 247 121
rect 407 297 465 309
rect 407 121 419 297
rect 453 121 465 297
rect 407 109 465 121
rect -465 -121 -407 -109
rect -465 -297 -453 -121
rect -419 -297 -407 -121
rect -465 -309 -407 -297
rect -247 -121 -189 -109
rect -247 -297 -235 -121
rect -201 -297 -189 -121
rect -247 -309 -189 -297
rect -29 -121 29 -109
rect -29 -297 -17 -121
rect 17 -297 29 -121
rect -29 -309 29 -297
rect 189 -121 247 -109
rect 189 -297 201 -121
rect 235 -297 247 -121
rect 189 -309 247 -297
rect 407 -121 465 -109
rect 407 -297 419 -121
rect 453 -297 465 -121
rect 407 -309 465 -297
<< ndiffc >>
rect -453 121 -419 297
rect -235 121 -201 297
rect -17 121 17 297
rect 201 121 235 297
rect 419 121 453 297
rect -453 -297 -419 -121
rect -235 -297 -201 -121
rect -17 -297 17 -121
rect 201 -297 235 -121
rect 419 -297 453 -121
<< poly >>
rect -407 381 -247 397
rect -407 347 -391 381
rect -263 347 -247 381
rect -407 309 -247 347
rect -189 381 -29 397
rect -189 347 -173 381
rect -45 347 -29 381
rect -189 309 -29 347
rect 29 381 189 397
rect 29 347 45 381
rect 173 347 189 381
rect 29 309 189 347
rect 247 381 407 397
rect 247 347 263 381
rect 391 347 407 381
rect 247 309 407 347
rect -407 71 -247 109
rect -407 37 -391 71
rect -263 37 -247 71
rect -407 21 -247 37
rect -189 71 -29 109
rect -189 37 -173 71
rect -45 37 -29 71
rect -189 21 -29 37
rect 29 71 189 109
rect 29 37 45 71
rect 173 37 189 71
rect 29 21 189 37
rect 247 71 407 109
rect 247 37 263 71
rect 391 37 407 71
rect 247 21 407 37
rect -407 -37 -247 -21
rect -407 -71 -391 -37
rect -263 -71 -247 -37
rect -407 -109 -247 -71
rect -189 -37 -29 -21
rect -189 -71 -173 -37
rect -45 -71 -29 -37
rect -189 -109 -29 -71
rect 29 -37 189 -21
rect 29 -71 45 -37
rect 173 -71 189 -37
rect 29 -109 189 -71
rect 247 -37 407 -21
rect 247 -71 263 -37
rect 391 -71 407 -37
rect 247 -109 407 -71
rect -407 -347 -247 -309
rect -407 -381 -391 -347
rect -263 -381 -247 -347
rect -407 -397 -247 -381
rect -189 -347 -29 -309
rect -189 -381 -173 -347
rect -45 -381 -29 -347
rect -189 -397 -29 -381
rect 29 -347 189 -309
rect 29 -381 45 -347
rect 173 -381 189 -347
rect 29 -397 189 -381
rect 247 -347 407 -309
rect 247 -381 263 -347
rect 391 -381 407 -347
rect 247 -397 407 -381
<< polycont >>
rect -391 347 -263 381
rect -173 347 -45 381
rect 45 347 173 381
rect 263 347 391 381
rect -391 37 -263 71
rect -173 37 -45 71
rect 45 37 173 71
rect 263 37 391 71
rect -391 -71 -263 -37
rect -173 -71 -45 -37
rect 45 -71 173 -37
rect 263 -71 391 -37
rect -391 -381 -263 -347
rect -173 -381 -45 -347
rect 45 -381 173 -347
rect 263 -381 391 -347
<< locali >>
rect -407 347 -391 381
rect -263 347 -247 381
rect -189 347 -173 381
rect -45 347 -29 381
rect 29 347 45 381
rect 173 347 189 381
rect 247 347 263 381
rect 391 347 407 381
rect -453 297 -419 313
rect -453 105 -419 121
rect -235 297 -201 313
rect -235 105 -201 121
rect -17 297 17 313
rect -17 105 17 121
rect 201 297 235 313
rect 201 105 235 121
rect 419 297 453 313
rect 419 105 453 121
rect -407 37 -391 71
rect -263 37 -247 71
rect -189 37 -173 71
rect -45 37 -29 71
rect 29 37 45 71
rect 173 37 189 71
rect 247 37 263 71
rect 391 37 407 71
rect -407 -71 -391 -37
rect -263 -71 -247 -37
rect -189 -71 -173 -37
rect -45 -71 -29 -37
rect 29 -71 45 -37
rect 173 -71 189 -37
rect 247 -71 263 -37
rect 391 -71 407 -37
rect -453 -121 -419 -105
rect -453 -313 -419 -297
rect -235 -121 -201 -105
rect -235 -313 -201 -297
rect -17 -121 17 -105
rect -17 -313 17 -297
rect 201 -121 235 -105
rect 201 -313 235 -297
rect 419 -121 453 -105
rect 419 -313 453 -297
rect -407 -381 -391 -347
rect -263 -381 -247 -347
rect -189 -381 -173 -347
rect -45 -381 -29 -347
rect 29 -381 45 -347
rect 173 -381 189 -347
rect 247 -381 263 -347
rect 391 -381 407 -347
<< viali >>
rect -372 347 -282 381
rect -154 347 -64 381
rect 64 347 154 381
rect 282 347 372 381
rect -453 121 -419 297
rect -235 121 -201 297
rect -17 121 17 297
rect 201 121 235 297
rect 419 121 453 297
rect -372 37 -282 71
rect -154 37 -64 71
rect 64 37 154 71
rect 282 37 372 71
rect -372 -71 -282 -37
rect -154 -71 -64 -37
rect 64 -71 154 -37
rect 282 -71 372 -37
rect -453 -297 -419 -121
rect -235 -297 -201 -121
rect -17 -297 17 -121
rect 201 -297 235 -121
rect 419 -297 453 -121
rect -372 -381 -282 -347
rect -154 -381 -64 -347
rect 64 -381 154 -347
rect 282 -381 372 -347
<< metal1 >>
rect -384 381 -270 387
rect -384 347 -372 381
rect -282 347 -270 381
rect -384 341 -270 347
rect -166 381 -52 387
rect -166 347 -154 381
rect -64 347 -52 381
rect -166 341 -52 347
rect 52 381 166 387
rect 52 347 64 381
rect 154 347 166 381
rect 52 341 166 347
rect 270 381 384 387
rect 270 347 282 381
rect 372 347 384 381
rect 270 341 384 347
rect -459 297 -413 309
rect -459 121 -453 297
rect -419 121 -413 297
rect -459 109 -413 121
rect -241 297 -195 309
rect -241 121 -235 297
rect -201 121 -195 297
rect -241 109 -195 121
rect -23 297 23 309
rect -23 121 -17 297
rect 17 121 23 297
rect -23 109 23 121
rect 195 297 241 309
rect 195 121 201 297
rect 235 121 241 297
rect 195 109 241 121
rect 413 297 459 309
rect 413 121 419 297
rect 453 121 459 297
rect 413 109 459 121
rect -384 71 -270 77
rect -384 37 -372 71
rect -282 37 -270 71
rect -384 31 -270 37
rect -166 71 -52 77
rect -166 37 -154 71
rect -64 37 -52 71
rect -166 31 -52 37
rect 52 71 166 77
rect 52 37 64 71
rect 154 37 166 71
rect 52 31 166 37
rect 270 71 384 77
rect 270 37 282 71
rect 372 37 384 71
rect 270 31 384 37
rect -384 -37 -270 -31
rect -384 -71 -372 -37
rect -282 -71 -270 -37
rect -384 -77 -270 -71
rect -166 -37 -52 -31
rect -166 -71 -154 -37
rect -64 -71 -52 -37
rect -166 -77 -52 -71
rect 52 -37 166 -31
rect 52 -71 64 -37
rect 154 -71 166 -37
rect 52 -77 166 -71
rect 270 -37 384 -31
rect 270 -71 282 -37
rect 372 -71 384 -37
rect 270 -77 384 -71
rect -459 -121 -413 -109
rect -459 -297 -453 -121
rect -419 -297 -413 -121
rect -459 -309 -413 -297
rect -241 -121 -195 -109
rect -241 -297 -235 -121
rect -201 -297 -195 -121
rect -241 -309 -195 -297
rect -23 -121 23 -109
rect -23 -297 -17 -121
rect 17 -297 23 -121
rect -23 -309 23 -297
rect 195 -121 241 -109
rect 195 -297 201 -121
rect 235 -297 241 -121
rect 195 -309 241 -297
rect 413 -121 459 -109
rect 413 -297 419 -121
rect 453 -297 459 -121
rect 413 -309 459 -297
rect -384 -347 -270 -341
rect -384 -381 -372 -347
rect -282 -381 -270 -347
rect -384 -387 -270 -381
rect -166 -347 -52 -341
rect -166 -381 -154 -347
rect -64 -381 -52 -347
rect -166 -387 -52 -381
rect 52 -347 166 -341
rect 52 -381 64 -347
rect 154 -381 166 -347
rect 52 -387 166 -381
rect 270 -347 384 -341
rect 270 -381 282 -347
rect 372 -381 384 -347
rect 270 -387 384 -381
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1 l 0.8 m 2 nf 4 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 70 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
