magic
tech sky130A
magscale 1 2
timestamp 1729224540
<< nmos >>
rect -578 55 -418 255
rect -246 55 -86 255
rect 86 55 246 255
rect 418 55 578 255
rect -578 -255 -418 -55
rect -246 -255 -86 -55
rect 86 -255 246 -55
rect 418 -255 578 -55
<< ndiff >>
rect -636 243 -578 255
rect -636 67 -624 243
rect -590 67 -578 243
rect -636 55 -578 67
rect -418 243 -360 255
rect -418 67 -406 243
rect -372 67 -360 243
rect -418 55 -360 67
rect -304 243 -246 255
rect -304 67 -292 243
rect -258 67 -246 243
rect -304 55 -246 67
rect -86 243 -28 255
rect -86 67 -74 243
rect -40 67 -28 243
rect -86 55 -28 67
rect 28 243 86 255
rect 28 67 40 243
rect 74 67 86 243
rect 28 55 86 67
rect 246 243 304 255
rect 246 67 258 243
rect 292 67 304 243
rect 246 55 304 67
rect 360 243 418 255
rect 360 67 372 243
rect 406 67 418 243
rect 360 55 418 67
rect 578 243 636 255
rect 578 67 590 243
rect 624 67 636 243
rect 578 55 636 67
rect -636 -67 -578 -55
rect -636 -243 -624 -67
rect -590 -243 -578 -67
rect -636 -255 -578 -243
rect -418 -67 -360 -55
rect -418 -243 -406 -67
rect -372 -243 -360 -67
rect -418 -255 -360 -243
rect -304 -67 -246 -55
rect -304 -243 -292 -67
rect -258 -243 -246 -67
rect -304 -255 -246 -243
rect -86 -67 -28 -55
rect -86 -243 -74 -67
rect -40 -243 -28 -67
rect -86 -255 -28 -243
rect 28 -67 86 -55
rect 28 -243 40 -67
rect 74 -243 86 -67
rect 28 -255 86 -243
rect 246 -67 304 -55
rect 246 -243 258 -67
rect 292 -243 304 -67
rect 246 -255 304 -243
rect 360 -67 418 -55
rect 360 -243 372 -67
rect 406 -243 418 -67
rect 360 -255 418 -243
rect 578 -67 636 -55
rect 578 -243 590 -67
rect 624 -243 636 -67
rect 578 -255 636 -243
<< ndiffc >>
rect -624 67 -590 243
rect -406 67 -372 243
rect -292 67 -258 243
rect -74 67 -40 243
rect 40 67 74 243
rect 258 67 292 243
rect 372 67 406 243
rect 590 67 624 243
rect -624 -243 -590 -67
rect -406 -243 -372 -67
rect -292 -243 -258 -67
rect -74 -243 -40 -67
rect 40 -243 74 -67
rect 258 -243 292 -67
rect 372 -243 406 -67
rect 590 -243 624 -67
<< poly >>
rect -578 327 -418 343
rect -578 293 -562 327
rect -434 293 -418 327
rect -578 255 -418 293
rect -246 327 -86 343
rect -246 293 -230 327
rect -102 293 -86 327
rect -246 255 -86 293
rect 86 327 246 343
rect 86 293 102 327
rect 230 293 246 327
rect 86 255 246 293
rect 418 327 578 343
rect 418 293 434 327
rect 562 293 578 327
rect 418 255 578 293
rect -578 17 -418 55
rect -578 -17 -562 17
rect -434 -17 -418 17
rect -578 -55 -418 -17
rect -246 17 -86 55
rect -246 -17 -230 17
rect -102 -17 -86 17
rect -246 -55 -86 -17
rect 86 17 246 55
rect 86 -17 102 17
rect 230 -17 246 17
rect 86 -55 246 -17
rect 418 17 578 55
rect 418 -17 434 17
rect 562 -17 578 17
rect 418 -55 578 -17
rect -578 -293 -418 -255
rect -578 -327 -562 -293
rect -434 -327 -418 -293
rect -578 -343 -418 -327
rect -246 -293 -86 -255
rect -246 -327 -230 -293
rect -102 -327 -86 -293
rect -246 -343 -86 -327
rect 86 -293 246 -255
rect 86 -327 102 -293
rect 230 -327 246 -293
rect 86 -343 246 -327
rect 418 -293 578 -255
rect 418 -327 434 -293
rect 562 -327 578 -293
rect 418 -343 578 -327
<< polycont >>
rect -562 293 -434 327
rect -230 293 -102 327
rect 102 293 230 327
rect 434 293 562 327
rect -562 -17 -434 17
rect -230 -17 -102 17
rect 102 -17 230 17
rect 434 -17 562 17
rect -562 -327 -434 -293
rect -230 -327 -102 -293
rect 102 -327 230 -293
rect 434 -327 562 -293
<< locali >>
rect -578 293 -562 327
rect -434 293 -418 327
rect -246 293 -230 327
rect -102 293 -86 327
rect 86 293 102 327
rect 230 293 246 327
rect 418 293 434 327
rect 562 293 578 327
rect -624 243 -590 259
rect -624 51 -590 67
rect -406 243 -372 259
rect -406 51 -372 67
rect -292 243 -258 259
rect -292 51 -258 67
rect -74 243 -40 259
rect -74 51 -40 67
rect 40 243 74 259
rect 40 51 74 67
rect 258 243 292 259
rect 258 51 292 67
rect 372 243 406 259
rect 372 51 406 67
rect 590 243 624 259
rect 590 51 624 67
rect -578 -17 -562 17
rect -434 -17 -418 17
rect -246 -17 -230 17
rect -102 -17 -86 17
rect 86 -17 102 17
rect 230 -17 246 17
rect 418 -17 434 17
rect 562 -17 578 17
rect -624 -67 -590 -51
rect -624 -259 -590 -243
rect -406 -67 -372 -51
rect -406 -259 -372 -243
rect -292 -67 -258 -51
rect -292 -259 -258 -243
rect -74 -67 -40 -51
rect -74 -259 -40 -243
rect 40 -67 74 -51
rect 40 -259 74 -243
rect 258 -67 292 -51
rect 258 -259 292 -243
rect 372 -67 406 -51
rect 372 -259 406 -243
rect 590 -67 624 -51
rect 590 -259 624 -243
rect -578 -327 -562 -293
rect -434 -327 -418 -293
rect -246 -327 -230 -293
rect -102 -327 -86 -293
rect 86 -327 102 -293
rect 230 -327 246 -293
rect 418 -327 434 -293
rect 562 -327 578 -293
<< viali >>
rect -543 293 -453 327
rect -211 293 -121 327
rect 121 293 211 327
rect 453 293 543 327
rect -624 67 -590 243
rect -406 67 -372 243
rect -292 67 -258 243
rect -74 67 -40 243
rect 40 67 74 243
rect 258 67 292 243
rect 372 67 406 243
rect 590 67 624 243
rect -543 -17 -453 17
rect -211 -17 -121 17
rect 121 -17 211 17
rect 453 -17 543 17
rect -624 -243 -590 -67
rect -406 -243 -372 -67
rect -292 -243 -258 -67
rect -74 -243 -40 -67
rect 40 -243 74 -67
rect 258 -243 292 -67
rect 372 -243 406 -67
rect 590 -243 624 -67
rect -543 -327 -453 -293
rect -211 -327 -121 -293
rect 121 -327 211 -293
rect 453 -327 543 -293
<< metal1 >>
rect -555 327 -441 333
rect -555 293 -543 327
rect -453 293 -441 327
rect -555 287 -441 293
rect -223 327 -109 333
rect -223 293 -211 327
rect -121 293 -109 327
rect -223 287 -109 293
rect 109 327 223 333
rect 109 293 121 327
rect 211 293 223 327
rect 109 287 223 293
rect 441 327 555 333
rect 441 293 453 327
rect 543 293 555 327
rect 441 287 555 293
rect -630 243 -584 255
rect -630 67 -624 243
rect -590 67 -584 243
rect -630 55 -584 67
rect -412 243 -366 255
rect -412 67 -406 243
rect -372 67 -366 243
rect -412 55 -366 67
rect -298 243 -252 255
rect -298 67 -292 243
rect -258 67 -252 243
rect -298 55 -252 67
rect -80 243 -34 255
rect -80 67 -74 243
rect -40 67 -34 243
rect -80 55 -34 67
rect 34 243 80 255
rect 34 67 40 243
rect 74 67 80 243
rect 34 55 80 67
rect 252 243 298 255
rect 252 67 258 243
rect 292 67 298 243
rect 252 55 298 67
rect 366 243 412 255
rect 366 67 372 243
rect 406 67 412 243
rect 366 55 412 67
rect 584 243 630 255
rect 584 67 590 243
rect 624 67 630 243
rect 584 55 630 67
rect -555 17 -441 23
rect -555 -17 -543 17
rect -453 -17 -441 17
rect -555 -23 -441 -17
rect -223 17 -109 23
rect -223 -17 -211 17
rect -121 -17 -109 17
rect -223 -23 -109 -17
rect 109 17 223 23
rect 109 -17 121 17
rect 211 -17 223 17
rect 109 -23 223 -17
rect 441 17 555 23
rect 441 -17 453 17
rect 543 -17 555 17
rect 441 -23 555 -17
rect -630 -67 -584 -55
rect -630 -243 -624 -67
rect -590 -243 -584 -67
rect -630 -255 -584 -243
rect -412 -67 -366 -55
rect -412 -243 -406 -67
rect -372 -243 -366 -67
rect -412 -255 -366 -243
rect -298 -67 -252 -55
rect -298 -243 -292 -67
rect -258 -243 -252 -67
rect -298 -255 -252 -243
rect -80 -67 -34 -55
rect -80 -243 -74 -67
rect -40 -243 -34 -67
rect -80 -255 -34 -243
rect 34 -67 80 -55
rect 34 -243 40 -67
rect 74 -243 80 -67
rect 34 -255 80 -243
rect 252 -67 298 -55
rect 252 -243 258 -67
rect 292 -243 298 -67
rect 252 -255 298 -243
rect 366 -67 412 -55
rect 366 -243 372 -67
rect 406 -243 412 -67
rect 366 -255 412 -243
rect 584 -67 630 -55
rect 584 -243 590 -67
rect 624 -243 630 -67
rect 584 -255 630 -243
rect -555 -293 -441 -287
rect -555 -327 -543 -293
rect -453 -327 -441 -293
rect -555 -333 -441 -327
rect -223 -293 -109 -287
rect -223 -327 -211 -293
rect -121 -327 -109 -293
rect -223 -333 -109 -327
rect 109 -293 223 -287
rect 109 -327 121 -293
rect 211 -327 223 -293
rect 109 -333 223 -327
rect 441 -293 555 -287
rect 441 -327 453 -293
rect 543 -327 555 -293
rect 441 -333 555 -327
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1 l 0.8 m 2 nf 4 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 1 doverlap 0 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 70 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
