magic
tech sky130A
magscale 1 2
timestamp 1729239931
<< error_p >>
rect -444 399 -372 405
rect -172 399 -100 405
rect 100 399 172 405
rect 372 399 444 405
rect -444 365 -432 399
rect -172 365 -160 399
rect 100 365 112 399
rect 372 365 384 399
rect -444 359 -372 365
rect -172 359 -100 365
rect 100 359 172 365
rect 372 359 444 365
rect -552 18 552 236
rect -444 -37 -372 -31
rect -172 -37 -100 -31
rect 100 -37 172 -31
rect 372 -37 444 -31
rect -444 -71 -432 -37
rect -172 -71 -160 -37
rect 100 -71 112 -37
rect 372 -71 384 -37
rect -444 -77 -372 -71
rect -172 -77 -100 -71
rect 100 -77 172 -71
rect 372 -77 444 -71
rect -444 -365 -372 -359
rect -172 -365 -100 -359
rect 100 -365 172 -359
rect 372 -365 444 -359
rect -444 -399 -432 -365
rect -172 -399 -160 -365
rect 100 -399 112 -365
rect 372 -399 384 -365
rect -444 -405 -372 -399
rect -172 -405 -100 -399
rect 100 -405 172 -399
rect 372 -405 444 -399
<< nwell >>
rect -552 18 552 418
rect -552 -418 552 -18
<< pmos >>
rect -458 118 -358 318
rect -186 118 -86 318
rect 86 118 186 318
rect 358 118 458 318
rect -458 -318 -358 -118
rect -186 -318 -86 -118
rect 86 -318 186 -118
rect 358 -318 458 -118
<< pdiff >>
rect -516 306 -458 318
rect -516 130 -504 306
rect -470 130 -458 306
rect -516 118 -458 130
rect -358 306 -300 318
rect -358 130 -346 306
rect -312 130 -300 306
rect -358 118 -300 130
rect -244 306 -186 318
rect -244 130 -232 306
rect -198 130 -186 306
rect -244 118 -186 130
rect -86 306 -28 318
rect -86 130 -74 306
rect -40 130 -28 306
rect -86 118 -28 130
rect 28 306 86 318
rect 28 130 40 306
rect 74 130 86 306
rect 28 118 86 130
rect 186 306 244 318
rect 186 130 198 306
rect 232 130 244 306
rect 186 118 244 130
rect 300 306 358 318
rect 300 130 312 306
rect 346 130 358 306
rect 300 118 358 130
rect 458 306 516 318
rect 458 130 470 306
rect 504 130 516 306
rect 458 118 516 130
rect -516 -130 -458 -118
rect -516 -306 -504 -130
rect -470 -306 -458 -130
rect -516 -318 -458 -306
rect -358 -130 -300 -118
rect -358 -306 -346 -130
rect -312 -306 -300 -130
rect -358 -318 -300 -306
rect -244 -130 -186 -118
rect -244 -306 -232 -130
rect -198 -306 -186 -130
rect -244 -318 -186 -306
rect -86 -130 -28 -118
rect -86 -306 -74 -130
rect -40 -306 -28 -130
rect -86 -318 -28 -306
rect 28 -130 86 -118
rect 28 -306 40 -130
rect 74 -306 86 -130
rect 28 -318 86 -306
rect 186 -130 244 -118
rect 186 -306 198 -130
rect 232 -306 244 -130
rect 186 -318 244 -306
rect 300 -130 358 -118
rect 300 -306 312 -130
rect 346 -306 358 -130
rect 300 -318 358 -306
rect 458 -130 516 -118
rect 458 -306 470 -130
rect 504 -306 516 -130
rect 458 -318 516 -306
<< pdiffc >>
rect -504 130 -470 306
rect -346 130 -312 306
rect -232 130 -198 306
rect -74 130 -40 306
rect 40 130 74 306
rect 198 130 232 306
rect 312 130 346 306
rect 470 130 504 306
rect -504 -306 -470 -130
rect -346 -306 -312 -130
rect -232 -306 -198 -130
rect -74 -306 -40 -130
rect 40 -306 74 -130
rect 198 -306 232 -130
rect 312 -306 346 -130
rect 470 -306 504 -130
<< poly >>
rect -458 399 -358 415
rect -458 365 -442 399
rect -374 365 -358 399
rect -458 318 -358 365
rect -186 399 -86 415
rect -186 365 -170 399
rect -102 365 -86 399
rect -186 318 -86 365
rect 86 399 186 415
rect 86 365 102 399
rect 170 365 186 399
rect 86 318 186 365
rect 358 399 458 415
rect 358 365 374 399
rect 442 365 458 399
rect 358 318 458 365
rect -458 71 -358 118
rect -458 37 -442 71
rect -374 37 -358 71
rect -458 21 -358 37
rect -186 71 -86 118
rect -186 37 -170 71
rect -102 37 -86 71
rect -186 21 -86 37
rect 86 71 186 118
rect 86 37 102 71
rect 170 37 186 71
rect 86 21 186 37
rect 358 71 458 118
rect 358 37 374 71
rect 442 37 458 71
rect 358 21 458 37
rect -458 -37 -358 -21
rect -458 -71 -442 -37
rect -374 -71 -358 -37
rect -458 -118 -358 -71
rect -186 -37 -86 -21
rect -186 -71 -170 -37
rect -102 -71 -86 -37
rect -186 -118 -86 -71
rect 86 -37 186 -21
rect 86 -71 102 -37
rect 170 -71 186 -37
rect 86 -118 186 -71
rect 358 -37 458 -21
rect 358 -71 374 -37
rect 442 -71 458 -37
rect 358 -118 458 -71
rect -458 -365 -358 -318
rect -458 -399 -442 -365
rect -374 -399 -358 -365
rect -458 -415 -358 -399
rect -186 -365 -86 -318
rect -186 -399 -170 -365
rect -102 -399 -86 -365
rect -186 -415 -86 -399
rect 86 -365 186 -318
rect 86 -399 102 -365
rect 170 -399 186 -365
rect 86 -415 186 -399
rect 358 -365 458 -318
rect 358 -399 374 -365
rect 442 -399 458 -365
rect 358 -415 458 -399
<< polycont >>
rect -442 365 -374 399
rect -170 365 -102 399
rect 102 365 170 399
rect 374 365 442 399
rect -442 37 -374 71
rect -170 37 -102 71
rect 102 37 170 71
rect 374 37 442 71
rect -442 -71 -374 -37
rect -170 -71 -102 -37
rect 102 -71 170 -37
rect 374 -71 442 -37
rect -442 -399 -374 -365
rect -170 -399 -102 -365
rect 102 -399 170 -365
rect 374 -399 442 -365
<< locali >>
rect -458 365 -442 399
rect -374 365 -358 399
rect -186 365 -170 399
rect -102 365 -86 399
rect 86 365 102 399
rect 170 365 186 399
rect 358 365 374 399
rect 442 365 458 399
rect -504 306 -470 322
rect -504 114 -470 130
rect -346 306 -312 322
rect -346 114 -312 130
rect -232 306 -198 322
rect -232 114 -198 130
rect -74 306 -40 322
rect -74 114 -40 130
rect 40 306 74 322
rect 40 114 74 130
rect 198 306 232 322
rect 198 114 232 130
rect 312 306 346 322
rect 312 114 346 130
rect 470 306 504 322
rect 470 114 504 130
rect -458 37 -442 71
rect -374 37 -358 71
rect -186 37 -170 71
rect -102 37 -86 71
rect 86 37 102 71
rect 170 37 186 71
rect 358 37 374 71
rect 442 37 458 71
rect -458 -71 -442 -37
rect -374 -71 -358 -37
rect -186 -71 -170 -37
rect -102 -71 -86 -37
rect 86 -71 102 -37
rect 170 -71 186 -37
rect 358 -71 374 -37
rect 442 -71 458 -37
rect -504 -130 -470 -114
rect -504 -322 -470 -306
rect -346 -130 -312 -114
rect -346 -322 -312 -306
rect -232 -130 -198 -114
rect -232 -322 -198 -306
rect -74 -130 -40 -114
rect -74 -322 -40 -306
rect 40 -130 74 -114
rect 40 -322 74 -306
rect 198 -130 232 -114
rect 198 -322 232 -306
rect 312 -130 346 -114
rect 312 -322 346 -306
rect 470 -130 504 -114
rect 470 -322 504 -306
rect -458 -399 -442 -365
rect -374 -399 -358 -365
rect -186 -399 -170 -365
rect -102 -399 -86 -365
rect 86 -399 102 -365
rect 170 -399 186 -365
rect 358 -399 374 -365
rect 442 -399 458 -365
<< viali >>
rect -432 365 -384 399
rect -160 365 -112 399
rect 112 365 160 399
rect 384 365 432 399
rect -504 130 -470 306
rect -346 130 -312 306
rect -232 130 -198 306
rect -74 130 -40 306
rect 40 130 74 306
rect 198 130 232 306
rect 312 130 346 306
rect 470 130 504 306
rect -432 37 -384 71
rect -160 37 -112 71
rect 112 37 160 71
rect 384 37 432 71
rect -432 -71 -384 -37
rect -160 -71 -112 -37
rect 112 -71 160 -37
rect 384 -71 432 -37
rect -504 -306 -470 -130
rect -346 -306 -312 -130
rect -232 -306 -198 -130
rect -74 -306 -40 -130
rect 40 -306 74 -130
rect 198 -306 232 -130
rect 312 -306 346 -130
rect 470 -306 504 -130
rect -432 -399 -384 -365
rect -160 -399 -112 -365
rect 112 -399 160 -365
rect 384 -399 432 -365
<< metal1 >>
rect -444 399 -372 405
rect -444 365 -432 399
rect -384 365 -372 399
rect -444 359 -372 365
rect -172 399 -100 405
rect -172 365 -160 399
rect -112 365 -100 399
rect -172 359 -100 365
rect 100 399 172 405
rect 100 365 112 399
rect 160 365 172 399
rect 100 359 172 365
rect 372 399 444 405
rect 372 365 384 399
rect 432 365 444 399
rect 372 359 444 365
rect -510 306 -464 318
rect -510 130 -504 306
rect -470 130 -464 306
rect -510 118 -464 130
rect -352 306 -306 318
rect -352 130 -346 306
rect -312 130 -306 306
rect -352 118 -306 130
rect -238 306 -192 318
rect -238 130 -232 306
rect -198 130 -192 306
rect -238 118 -192 130
rect -80 306 -34 318
rect -80 130 -74 306
rect -40 130 -34 306
rect -80 118 -34 130
rect 34 306 80 318
rect 34 130 40 306
rect 74 130 80 306
rect 34 118 80 130
rect 192 306 238 318
rect 192 130 198 306
rect 232 130 238 306
rect 192 118 238 130
rect 306 306 352 318
rect 306 130 312 306
rect 346 130 352 306
rect 306 118 352 130
rect 464 306 510 318
rect 464 130 470 306
rect 504 130 510 306
rect 464 118 510 130
rect -444 71 -372 77
rect -444 37 -432 71
rect -384 37 -372 71
rect -444 31 -372 37
rect -172 71 -100 77
rect -172 37 -160 71
rect -112 37 -100 71
rect -172 31 -100 37
rect 100 71 172 77
rect 100 37 112 71
rect 160 37 172 71
rect 100 31 172 37
rect 372 71 444 77
rect 372 37 384 71
rect 432 37 444 71
rect 372 31 444 37
rect -444 -37 -372 -31
rect -444 -71 -432 -37
rect -384 -71 -372 -37
rect -444 -77 -372 -71
rect -172 -37 -100 -31
rect -172 -71 -160 -37
rect -112 -71 -100 -37
rect -172 -77 -100 -71
rect 100 -37 172 -31
rect 100 -71 112 -37
rect 160 -71 172 -37
rect 100 -77 172 -71
rect 372 -37 444 -31
rect 372 -71 384 -37
rect 432 -71 444 -37
rect 372 -77 444 -71
rect -510 -130 -464 -118
rect -510 -306 -504 -130
rect -470 -306 -464 -130
rect -510 -318 -464 -306
rect -352 -130 -306 -118
rect -352 -306 -346 -130
rect -312 -306 -306 -130
rect -352 -318 -306 -306
rect -238 -130 -192 -118
rect -238 -306 -232 -130
rect -198 -306 -192 -130
rect -238 -318 -192 -306
rect -80 -130 -34 -118
rect -80 -306 -74 -130
rect -40 -306 -34 -130
rect -80 -318 -34 -306
rect 34 -130 80 -118
rect 34 -306 40 -130
rect 74 -306 80 -130
rect 34 -318 80 -306
rect 192 -130 238 -118
rect 192 -306 198 -130
rect 232 -306 238 -130
rect 192 -318 238 -306
rect 306 -130 352 -118
rect 306 -306 312 -130
rect 346 -306 352 -130
rect 306 -318 352 -306
rect 464 -130 510 -118
rect 464 -306 470 -130
rect 504 -306 510 -130
rect 464 -318 510 -306
rect -444 -365 -372 -359
rect -444 -399 -432 -365
rect -384 -399 -372 -365
rect -444 -405 -372 -399
rect -172 -365 -100 -359
rect -172 -399 -160 -365
rect -112 -399 -100 -365
rect -172 -405 -100 -399
rect 100 -365 172 -359
rect 100 -399 112 -365
rect 160 -399 172 -365
rect 100 -405 172 -399
rect 372 -365 444 -359
rect 372 -399 384 -365
rect 432 -399 444 -365
rect 372 -405 444 -399
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1 l 0.5 m 2 nf 4 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 0 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 70 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
